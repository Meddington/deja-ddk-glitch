library verilog;
use verilog.vl_types.all;
entity glitch_power_tb is
end glitch_power_tb;
